library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity ROM_OBJ_0 is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(10 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of ROM_OBJ_0 is
	type rom is array(0 to  2047) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"38",X"7C",X"C1",X"81",X"85",X"7C",X"38",X"00",X"01",X"01",X"FD",X"FD",X"41",X"01",X"00",X"00",
		X"61",X"F1",X"B9",X"99",X"9D",X"CD",X"45",X"00",X"8C",X"DD",X"F1",X"B1",X"91",X"85",X"04",X"00",
		X"08",X"FD",X"FD",X"C8",X"68",X"38",X"18",X"00",X"1C",X"BD",X"A1",X"A1",X"A1",X"E5",X"E4",X"00",
		X"0C",X"9D",X"91",X"91",X"D1",X"7D",X"3C",X"00",X"C0",X"E0",X"B0",X"9D",X"8D",X"C0",X"C0",X"00",
		X"0C",X"6D",X"99",X"99",X"B1",X"F1",X"6C",X"00",X"78",X"FC",X"95",X"91",X"91",X"F1",X"60",X"00",
		X"3D",X"7D",X"C8",X"88",X"C8",X"7D",X"3D",X"00",X"6C",X"FD",X"91",X"91",X"91",X"FD",X"FD",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"3D",X"7D",X"C8",X"88",X"C8",X"7D",X"3D",X"00",
		X"6C",X"FD",X"91",X"91",X"91",X"FD",X"FD",X"00",X"44",X"C5",X"81",X"81",X"C5",X"7C",X"38",X"00",
		X"38",X"7C",X"C5",X"81",X"81",X"FD",X"FD",X"00",X"81",X"91",X"91",X"91",X"FD",X"FD",X"00",X"00",
		X"80",X"90",X"90",X"90",X"90",X"FD",X"FD",X"00",X"9D",X"9D",X"91",X"81",X"C5",X"7C",X"38",X"00",
		X"FD",X"FD",X"10",X"10",X"10",X"FD",X"FD",X"00",X"81",X"81",X"FD",X"FD",X"81",X"81",X"00",X"00",
		X"FC",X"FD",X"01",X"01",X"01",X"05",X"04",X"00",X"81",X"C5",X"6D",X"3C",X"18",X"FD",X"FD",X"00",
		X"01",X"01",X"01",X"01",X"FD",X"FD",X"00",X"00",X"FD",X"FD",X"70",X"38",X"70",X"FD",X"FD",X"00",
		X"FD",X"FD",X"1C",X"38",X"70",X"FD",X"FD",X"00",X"7C",X"FD",X"81",X"81",X"81",X"FD",X"7C",X"00",
		X"70",X"F8",X"88",X"88",X"88",X"FD",X"FD",X"00",X"79",X"FC",X"8D",X"89",X"81",X"FD",X"7C",X"00",
		X"71",X"F5",X"9D",X"8C",X"88",X"FD",X"FD",X"00",X"0C",X"5D",X"D1",X"91",X"91",X"F5",X"64",X"00",
		X"80",X"80",X"FD",X"FD",X"80",X"80",X"00",X"00",X"FC",X"FD",X"01",X"01",X"01",X"FD",X"FC",X"00",
		X"F0",X"F8",X"1C",X"0D",X"1C",X"F8",X"F0",X"00",X"F8",X"FD",X"1C",X"38",X"1C",X"FD",X"F8",X"00",
		X"C5",X"ED",X"7C",X"38",X"7C",X"ED",X"C5",X"00",X"C0",X"F0",X"1D",X"1D",X"F0",X"C0",X"00",X"00",
		X"C1",X"E1",X"F1",X"B9",X"9D",X"8D",X"85",X"00",X"10",X"10",X"10",X"10",X"10",X"10",X"10",X"00",
		X"00",X"00",X"00",X"00",X"08",X"0C",X"0D",X"0F",X"00",X"00",X"80",X"00",X"08",X"18",X"38",X"78",
		X"07",X"02",X"02",X"00",X"00",X"00",X"00",X"00",X"70",X"40",X"C0",X"80",X"80",X"00",X"00",X"00",
		X"04",X"0F",X"0F",X"0F",X"0F",X"0F",X"07",X"07",X"20",X"F0",X"F0",X"F0",X"F0",X"F0",X"E0",X"E0",
		X"0F",X"0F",X"0F",X"0F",X"0F",X"0E",X"07",X"00",X"F0",X"F0",X"F0",X"F0",X"F0",X"B0",X"E0",X"00",
		X"00",X"00",X"00",X"00",X"04",X"0C",X"00",X"00",X"00",X"00",X"80",X"00",X"10",X"58",X"20",X"10",
		X"00",X"00",X"00",X"0C",X"04",X"02",X"00",X"00",X"10",X"10",X"20",X"18",X"10",X"C0",X"80",X"00",
		X"00",X"02",X"00",X"08",X"18",X"0C",X"00",X"00",X"00",X"00",X"80",X"08",X"0C",X"58",X"20",X"10",
		X"00",X"00",X"00",X"0C",X"18",X"0A",X"02",X"00",X"10",X"10",X"20",X"18",X"0C",X"C8",X"C0",X"80",
		X"00",X"00",X"00",X"08",X"18",X"0C",X"00",X"00",X"00",X"40",X"80",X"08",X"0C",X"58",X"20",X"10",
		X"00",X"08",X"18",X"0C",X"00",X"02",X"02",X"00",X"10",X"18",X"2C",X"18",X"00",X"C0",X"C0",X"80",
		X"7E",X"D7",X"B3",X"F7",X"5F",X"CC",X"D8",X"F8",X"FB",X"DA",X"9B",X"BF",X"FF",X"41",X"00",X"00",
		X"E8",X"B8",X"98",X"BC",X"F8",X"10",X"00",X"00",X"B8",X"9C",X"B8",X"F8",X"58",X"C8",X"DC",X"F8",
		X"78",X"F8",X"DC",X"97",X"B3",X"F7",X"DF",X"76",X"00",X"00",X"41",X"FF",X"F7",X"B3",X"97",X"BD",
		X"00",X"00",X"10",X"F8",X"BD",X"98",X"B8",X"E8",X"77",X"FE",X"BC",X"FE",X"EF",X"E7",X"EE",X"7F",
		X"00",X"10",X"38",X"10",X"01",X"07",X"01",X"17",X"00",X"00",X"20",X"70",X"20",X"00",X"08",X"AC",
		X"3A",X"10",X"00",X"02",X"13",X"3A",X"10",X"00",X"C8",X"80",X"04",X"0D",X"84",X"12",X"38",X"10",
		X"00",X"1C",X"3D",X"1D",X"3D",X"1C",X"00",X"00",X"67",X"3C",X"3C",X"7C",X"3C",X"3C",X"67",X"00",
		X"3C",X"41",X"82",X"A6",X"A6",X"9A",X"41",X"3C",X"FF",X"82",X"82",X"82",X"82",X"82",X"82",X"FF",
		X"01",X"03",X"05",X"0F",X"05",X"07",X"05",X"07",X"40",X"C0",X"60",X"F0",X"60",X"E0",X"60",X"E0",
		X"07",X"07",X"07",X"0F",X"07",X"07",X"03",X"02",X"E0",X"E0",X"E0",X"F0",X"E0",X"E0",X"C0",X"80",
		X"02",X"02",X"00",X"00",X"00",X"08",X"00",X"00",X"38",X"38",X"38",X"38",X"D0",X"18",X"18",X"18",
		X"04",X"04",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"90",X"80",X"00",X"00",X"00",X"00",X"00",
		X"00",X"01",X"00",X"00",X"00",X"04",X"04",X"00",X"38",X"18",X"18",X"58",X"50",X"58",X"18",X"38",
		X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"08",X"38",X"38",X"38",X"38",X"30",X"B8",X"38",X"38",
		X"00",X"00",X"00",X"03",X"0D",X"18",X"18",X"18",X"00",X"00",X"00",X"C0",X"70",X"18",X"C8",X"00",
		X"0D",X"02",X"00",X"08",X"00",X"00",X"00",X"00",X"78",X"F8",X"78",X"30",X"78",X"78",X"38",X"38",
		X"07",X"08",X"08",X"08",X"07",X"00",X"07",X"08",X"C0",X"20",X"20",X"20",X"C0",X"00",X"C0",X"20",
		X"08",X"08",X"07",X"00",X"00",X"0F",X"04",X"00",X"20",X"20",X"C0",X"00",X"20",X"E0",X"20",X"00",
		X"07",X"08",X"08",X"07",X"00",X"07",X"08",X"08",X"C0",X"20",X"20",X"C0",X"00",X"C0",X"20",X"20",
		X"07",X"00",X"05",X"0A",X"08",X"08",X"04",X"00",X"C0",X"00",X"20",X"20",X"A0",X"60",X"20",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"20",X"20",X"20",X"20",X"21",X"26",X"22",
		X"00",X"00",X"00",X"00",X"03",X"03",X"00",X"00",X"40",X"41",X"06",X"02",X"02",X"02",X"42",X"20",
		X"02",X"03",X"62",X"90",X"97",X"7F",X"3B",X"3E",X"E0",X"FA",X"FB",X"FF",X"FD",X"FF",X"FC",X"E4",
		X"3E",X"3B",X"7F",X"97",X"90",X"62",X"03",X"02",X"E4",X"E4",X"FF",X"FD",X"FF",X"FB",X"FA",X"E0",
		X"00",X"00",X"10",X"3C",X"01",X"07",X"1F",X"1F",X"00",X"00",X"04",X"1D",X"30",X"E0",X"E0",X"E0",
		X"1F",X"1F",X"07",X"01",X"3C",X"10",X"00",X"00",X"E0",X"E0",X"E0",X"30",X"1D",X"04",X"00",X"00",
		X"00",X"00",X"00",X"10",X"3D",X"07",X"1F",X"1F",X"00",X"00",X"00",X"10",X"38",X"EC",X"E3",X"E0",
		X"1F",X"1F",X"07",X"3D",X"10",X"00",X"00",X"00",X"E0",X"E3",X"EC",X"38",X"10",X"00",X"00",X"00",
		X"00",X"00",X"08",X"1D",X"01",X"07",X"1F",X"1F",X"00",X"00",X"20",X"F0",X"80",X"C0",X"E0",X"E0",
		X"1F",X"1F",X"07",X"01",X"1D",X"08",X"00",X"00",X"E0",X"E0",X"C0",X"80",X"F0",X"20",X"00",X"00",
		X"00",X"10",X"30",X"10",X"18",X"0F",X"07",X"07",X"00",X"08",X"0C",X"08",X"18",X"F0",X"E0",X"E0",
		X"07",X"0F",X"17",X"13",X"33",X"10",X"00",X"00",X"E0",X"F0",X"E8",X"C8",X"CC",X"08",X"00",X"00",
		X"00",X"01",X"05",X"0C",X"18",X"0F",X"07",X"07",X"00",X"40",X"60",X"30",X"18",X"F0",X"E0",X"E0",
		X"07",X"0F",X"0F",X"0B",X"1B",X"08",X"00",X"00",X"E0",X"F0",X"F0",X"D0",X"D8",X"10",X"00",X"00",
		X"00",X"00",X"00",X"00",X"10",X"33",X"17",X"1F",X"00",X"00",X"00",X"00",X"08",X"CC",X"E8",X"F8",
		X"07",X"1F",X"17",X"33",X"13",X"00",X"00",X"00",X"E0",X"F8",X"E8",X"CC",X"C8",X"00",X"00",X"00",
		X"00",X"00",X"01",X"08",X"12",X"07",X"27",X"0F",X"00",X"00",X"40",X"10",X"88",X"E0",X"E4",X"F0",
		X"0F",X"27",X"07",X"12",X"08",X"01",X"00",X"00",X"F0",X"E4",X"E0",X"88",X"10",X"40",X"00",X"00",
		X"00",X"02",X"14",X"20",X"02",X"46",X"03",X"4F",X"00",X"80",X"28",X"04",X"80",X"A1",X"C0",X"F1",
		X"4F",X"03",X"46",X"02",X"20",X"14",X"02",X"00",X"F1",X"C0",X"A1",X"80",X"04",X"28",X"80",X"00",
		X"01",X"00",X"20",X"00",X"01",X"00",X"88",X"02",X"40",X"00",X"04",X"00",X"40",X"00",X"12",X"80",
		X"02",X"88",X"00",X"01",X"00",X"20",X"00",X"01",X"80",X"12",X"00",X"40",X"00",X"04",X"00",X"40",
		X"00",X"00",X"00",X"04",X"0A",X"03",X"07",X"07",X"00",X"00",X"00",X"10",X"88",X"C0",X"E0",X"E0",
		X"07",X"07",X"03",X"12",X"08",X"00",X"00",X"00",X"E0",X"E0",X"C0",X"88",X"10",X"00",X"00",X"00",
		X"00",X"02",X"00",X"00",X"00",X"01",X"04",X"22",X"00",X"80",X"00",X"00",X"00",X"20",X"90",X"C1",
		X"22",X"02",X"04",X"01",X"00",X"00",X"02",X"00",X"C1",X"C0",X"90",X"20",X"00",X"00",X"80",X"00",
		X"02",X"00",X"00",X"01",X"01",X"00",X"00",X"00",X"00",X"08",X"14",X"01",X"21",X"29",X"48",X"48",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"08",X"00",X"04",X"04",X"06",X"02",X"0A",X"08",
		X"02",X"03",X"07",X"07",X"0F",X"07",X"07",X"07",X"80",X"C0",X"E0",X"E0",X"F0",X"E0",X"E0",X"E0",
		X"07",X"05",X"05",X"05",X"0F",X"05",X"05",X"01",X"E0",X"60",X"E0",X"60",X"F0",X"60",X"E0",X"40",
		X"00",X"29",X"29",X"3F",X"08",X"08",X"0F",X"07",X"00",X"54",X"54",X"FC",X"10",X"10",X"F0",X"E0",
		X"07",X"3F",X"07",X"37",X"07",X"3F",X"03",X"00",X"EC",X"F0",X"EC",X"E0",X"EC",X"F0",X"CC",X"00",
		X"0F",X"1F",X"1F",X"1F",X"1F",X"0F",X"00",X"1F",X"F0",X"F0",X"F8",X"F8",X"F8",X"F0",X"00",X"F8",
		X"1F",X"1F",X"0F",X"07",X"00",X"00",X"00",X"00",X"F8",X"F8",X"F0",X"E0",X"00",X"00",X"00",X"00",
		X"00",X"00",X"0F",X"1F",X"1F",X"1F",X"0F",X"0F",X"00",X"00",X"F0",X"F8",X"F8",X"F8",X"F0",X"F0",
		X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"20",X"08",X"00",X"10",X"00",X"40",X"00",X"00",
		X"00",X"00",X"21",X"02",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"40",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"00",X"00",X"08",X"00",X"00",X"10",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"40",X"00",X"00",X"40",X"00",X"10",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"20",X"00",X"00",X"10",X"00",X"20",X"00",
		X"00",X"00",X"00",X"08",X"00",X"00",X"00",X"00",X"80",X"00",X"00",X"80",X"80",X"80",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"20",X"00",X"00",X"00",X"40",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"00",X"00",X"40",X"00",X"00",X"20",X"08",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"00",X"20",X"00",X"00",X"10",X"00",X"08",
		X"00",X"00",X"00",X"00",X"02",X"00",X"00",X"00",X"00",X"20",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"00",X"00",X"40",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"08",X"00",X"00",X"10",X"00",X"20",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"02",X"66",X"06",X"04",X"44",X"10",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"21",X"81",X"09",X"49",X"09",X"08",X"10",X"10",
		X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"02",X"02",X"84",X"04",X"00",X"21",X"46",X"02",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"86",X"02",X"0A",X"0A",X"40",X"44",X"14",X"14",
		X"00",X"00",X"00",X"00",X"18",X"00",X"0C",X"00",X"00",X"00",X"20",X"00",X"20",X"01",X"46",X"02",
		X"03",X"00",X"00",X"00",X"05",X"05",X"00",X"00",X"60",X"01",X"06",X"02",X"02",X"C2",X"82",X"20",
		X"C0",X"E0",X"E3",X"E3",X"E3",X"E3",X"E3",X"E3",X"00",X"00",X"00",X"80",X"80",X"80",X"80",X"80",
		X"E3",X"E3",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"80",X"80",X"FC",X"FD",X"FD",X"FD",X"01",X"00",
		X"7F",X"7F",X"FF",X"FF",X"C3",X"E3",X"E0",X"E0",X"0C",X"8D",X"BD",X"BD",X"FD",X"FD",X"F1",X"F8",
		X"E0",X"E0",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"F8",X"F8",X"FC",X"FD",X"FD",X"FD",X"01",X"00",
		X"3F",X"3F",X"FF",X"FF",X"C0",X"E0",X"E0",X"E0",X"F0",X"F8",X"FC",X"FD",X"0D",X"0D",X"0D",X"0D",
		X"E0",X"E0",X"FF",X"FF",X"3F",X"3F",X"00",X"00",X"0D",X"0D",X"FD",X"FD",X"F1",X"F8",X"08",X"00",
		X"00",X"00",X"08",X"40",X"48",X"00",X"00",X"00",X"00",X"08",X"04",X"31",X"29",X"49",X"28",X"0A",
		X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"02",X"2A",X"02",X"16",X"14",X"14",X"14",X"04",X"20",
		X"00",X"00",X"10",X"3B",X"7F",X"33",X"13",X"1F",X"00",X"00",X"08",X"DC",X"FD",X"FC",X"F8",X"F8",
		X"1F",X"13",X"33",X"7F",X"3B",X"10",X"00",X"00",X"F8",X"FC",X"FD",X"DC",X"08",X"00",X"00",X"00",
		X"00",X"30",X"77",X"7F",X"33",X"37",X"7F",X"7F",X"00",X"18",X"D8",X"FC",X"FC",X"F8",X"F8",X"F8",
		X"7F",X"7F",X"37",X"33",X"7F",X"77",X"30",X"00",X"F8",X"F8",X"F8",X"FC",X"FC",X"D8",X"18",X"00",
		X"30",X"63",X"FF",X"F8",X"BC",X"7F",X"7F",X"7F",X"0C",X"CC",X"FF",X"FF",X"FE",X"FD",X"FD",X"FD",
		X"7F",X"7F",X"7F",X"BC",X"F8",X"FF",X"63",X"30",X"FD",X"FD",X"FD",X"FE",X"FF",X"FF",X"CC",X"00",
		X"0C",X"0C",X"01",X"3A",X"68",X"DC",X"FD",X"FD",X"00",X"00",X"00",X"03",X"83",X"44",X"28",X"10",
		X"FD",X"DC",X"68",X"3A",X"01",X"0C",X"0C",X"00",X"28",X"44",X"83",X"03",X"00",X"00",X"00",X"00",
		X"C3",X"E3",X"E3",X"E3",X"E3",X"E3",X"E0",X"E0",X"FC",X"FD",X"FD",X"FD",X"0D",X"8D",X"8D",X"0D",
		X"F0",X"F8",X"3F",X"3F",X"0F",X"0F",X"00",X"00",X"3D",X"3D",X"F1",X"F8",X"C8",X"E0",X"20",X"00",
		X"C0",X"E0",X"E3",X"E3",X"E3",X"E3",X"E3",X"E3",X"0C",X"0D",X"0D",X"8D",X"8D",X"8D",X"8D",X"8D",
		X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"FD",X"FD",X"FD",X"FD",X"01",X"00",X"00",X"00",
		X"02",X"03",X"62",X"90",X"97",X"7F",X"3A",X"38",X"E0",X"FA",X"FB",X"FF",X"FD",X"FF",X"FC",X"E4",
		X"38",X"3A",X"7F",X"97",X"90",X"62",X"03",X"02",X"E4",X"E4",X"FF",X"FD",X"FF",X"FB",X"FA",X"E0");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
